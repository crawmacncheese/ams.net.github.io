*SPICE Netlist for circuit 0
C1 0 5 1nF
M1 1 4 0 0 NMOS W=1u L=1u
M2 2 2 6 6 PMOS W=1u L=1u
M3 5 3 6 6 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

