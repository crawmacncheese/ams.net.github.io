*SPICE Netlist for circuit 1
C1 2 5 1nF
C2 8 0 1nF
M1 4 10 0 0 NMOS W=1u L=1u
M2 11 11 12 12 PMOS W=1u L=1u
M3 2 6 12 12 PMOS W=1u L=1u
M4 7 8 3 3 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

