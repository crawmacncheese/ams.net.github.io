*SPICE Netlist for circuit 2
I1 13 0 DC 1mA
M3 5 14 0 0 NMOS W=1u L=1u
M4 3 15 0 0 NMOS W=1u L=1u
M7 1 1 12 12 PMOS W=1u L=1u
M8 3 1 16 16 PMOS W=1u L=1u
M1 1 2 2 2 NMOS W=1u L=1u
M2 4 7 2 2 NMOS W=1u L=1u
M6 5 4 16 16 PMOS W=1u L=1u
M5 4 4 11 11 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

