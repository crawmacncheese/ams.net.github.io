*SPICE Netlist for circuit 1


.OP
.END

