*SPICE Netlist for circuit 1
M7 18 4 0 0 NMOS W=1u L=1u
M2 19 20 0 0 NMOS W=1u L=1u
M3 21 9 0 0 NMOS W=1u L=1u
M10 5 1 15 15 PMOS W=1u L=1u
M4 17 12 2 2 NMOS W=1u L=1u
M1 7 2 2 2 NMOS W=1u L=1u
M5 5 3 19 19 NMOS W=1u L=1u
M9 7 6 22 22 PMOS W=1u L=1u
M11 8 23 7 7 PMOS W=1u L=1u
M6 8 24 21 21 NMOS W=1u L=1u
M8 17 22 22 22 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

