*SPICE Netlist for circuit 0
C1 1 5 1nF
C2 5 0 1nF
I1 2 0 DC 1mA
M2 3 7 2 2 NMOS W=1u L=1u
M1 1 5 2 2 NMOS W=1u L=1u
M3 3 3 9 9 PMOS W=1u L=1u
M4 1 8 9 9 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

