*SPICE Netlist for circuit 1
M1 5 5 6 6 PMOS W=1u L=1u
M3 6 2 7 7 PMOS W=1u L=1u
M2 8 3 7 7 PMOS W=1u L=1u
M4 1 4 8 8 PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

