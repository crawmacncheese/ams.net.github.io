*SPICE Netlist for circuit 0
M1 1 2 6 6 PMOS W=1u L=1u
M2 4 17 7 7 PMOS W=1u L=1u
M7 8 18 9 9 PMOS W=1u L=1u
M3 10 19 11 11 PMOS W=1u L=1u
M6 12 1 19 19 PMOS W=1u L=1u
M4 13 20 14 14 PMOS W=1u L=1u
M5 15 17 3 3 PMOS W=1u L=1u
M8 16 21 22 22 PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

