*SPICE Netlist for circuit 1
M1 4 4 5 5 PMOS W=1u L=1u
M2 5 2 6 6 PMOS W=1u L=1u
M3 1 3 6 6 PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

