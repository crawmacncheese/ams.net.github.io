*SPICE Netlist for circuit 1
M1 1 4 2 2 PMOS W=1u L=1u
M2 4 13 14 14 PMOS W=1u L=1u
M7 6 13 7 7 PMOS W=1u L=1u
M3 8 15 16 16 PMOS W=1u L=1u
M6 9 1 15 15 PMOS W=1u L=1u
M4 10 5 16 16 PMOS W=1u L=1u
M5 3 14 11 11 PMOS W=1u L=1u
M8 17 18 12 12 PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

