*SPICE Netlist for circuit 1
M7 3 5 0 0 NMOS W=1u L=1u
M2 20 21 0 0 NMOS W=1u L=1u
M3 22 6 0 0 NMOS W=1u L=1u
M9 8 1 23 23 PMOS W=1u L=1u
M10 7 2 15 15 PMOS W=1u L=1u
M4 18 12 3 3 NMOS W=1u L=1u
M1 8 13 3 3 NMOS W=1u L=1u
M5 7 4 20 20 NMOS W=1u L=1u
M11 9 24 8 8 PMOS W=1u L=1u
M6 9 25 22 22 NMOS W=1u L=1u
M8 17 23 23 23 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

