*SPICE Netlist for circuit 2


.OP
.END

