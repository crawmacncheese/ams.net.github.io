*SPICE Netlist for circuit 2
I1 14 0 DC 1mA
M3 6 3 0 0 NMOS W=1u L=1u
M4 4 15 0 0 NMOS W=1u L=1u
M7 1 1 13 13 PMOS W=1u L=1u
M8 4 1 16 16 PMOS W=1u L=1u
M1 1 2 2 2 NMOS W=1u L=1u
M2 5 8 2 2 NMOS W=1u L=1u
M6 6 5 16 16 PMOS W=1u L=1u
M5 5 5 12 12 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

